-- jtag_uart_8kw.vhd

-- Generated using ACDS version 17.0 595

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity jtag_uart_8kw is
	port (
		av_chipselect  : in  std_logic                     := '0';             -- av_avalon_jtag_slave.chipselect
		av_address     : in  std_logic                     := '0';             --                              .address
		av_read_n      : in  std_logic                     := '0';             --                              .read_n
		av_readdata    : out std_logic_vector(31 downto 0);                    --                              .readdata
		av_write_n     : in  std_logic                     := '0';             --                              .write_n
		av_writedata   : in  std_logic_vector(31 downto 0) := (others => '0'); --                              .writedata
		av_waitrequest : out std_logic;                                        --                              .waitrequest
		clk_clk                       : in  std_logic                     := '0';             --               av_clk.clk
		irq_irq                       : out std_logic;                                        --               av_irq.irq
		reset_reset_n                 : in  std_logic                     := '0'              --             av_reset.reset_n
	);
end entity jtag_uart_8kw;

architecture rtl of jtag_uart_8kw is
	component jtag_uart_8kw_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component jtag_uart_8kw_jtag_uart_0;

begin

	jtag_uart_0 : component jtag_uart_8kw_jtag_uart_0
		port map (
			clk            => clk_clk,                       --               clk.clk
			rst_n          => reset_reset_n,                 --             reset.reset_n
			av_chipselect  => av_chipselect,  -- avalon_jtag_slave.chipselect
			av_address     => av_address,     --                  .address
			av_read_n      => av_read_n,      --                  .read_n
			av_readdata    => av_readdata,    --                  .readdata
			av_write_n     => av_write_n,     --                  .write_n
			av_writedata   => av_writedata,   --                  .writedata
			av_waitrequest => av_waitrequest, --                  .waitrequest
			av_irq         => irq_irq                        --               irq.irq
		);

end architecture rtl; -- of jtag_uart_8kw
